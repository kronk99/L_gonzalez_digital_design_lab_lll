//Este archivo es el que controla el juego como tal. Instancia los módulos e interpreta el input del usuario

module Battleship();



endmodule